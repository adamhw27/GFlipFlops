module RegMux(r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15, sel, out);
	input [15:0] r0, r1, r2, r3, r4, r5, r6, r7, r8, r9, r10, r11, r12, r13, r14, r15;
	input [3:0] sel;
	output reg [15:0] out;

	always @(*) begin
	
		casex (sel)
		
		16'd0: 
			begin
			out = r0;
			end
			
		16'd1: 
			begin
			out = r1;
			end
			
		16'd2: 
			begin
			out = r2;
			end
			
		16'd3: 
			begin
			out = r3;
			end
			
		16'd4: 
			begin
			out = r4;
			end
			
		16'd5: 
			begin
			out = r5;
			end
			
		16'd6: 
			begin
			out = r6;
			end
			
		16'd7: 
			begin
			out = r7;
			end
			
		16'd8: 
			begin
			out = r8;
			end
			
		16'd9: 
			begin
			out = r9;
			end
			
		16'd10: 
			begin
			out = r10;
			end
			
		16'd11: 
			begin
			out = r11;
			end
			
		16'd12: 
			begin
			out = r12;
			end
			
		16'd13: 
			begin
			out = r13;
			end
			
		16'd14: 
			begin
			out = r14;
			end
			
		16'd15: 
			begin
			out = r15;
			end
		default:
			begin
			out = 16'd0;
			end
		
		endcase
			
	end
	
endmodule
	
		