module TwoInputMux(i0, i1, sel, out);
	input [15:0] i0, i1;
	input sel;
	output reg[15:0] out;
	
	
	always @* begin
		
		case (sel)
			16'd0:
				begin
				out <= i0;
				end
			16'd1:
				begin
				out <= i1;
				end
			default:
				begin
				out = 16'd0;
				end
		endcase
	end
endmodule